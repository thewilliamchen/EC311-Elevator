`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:58:51 11/29/2016 
// Design Name: 
// Module Name:    register_3b 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

//use the mux to feed into this, mux toggles switch/btn
module register_3b(
    input [2:0] in,
	 input clock,
    output [2:0] out
    );


endmodule
